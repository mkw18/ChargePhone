library verilog;
use verilog.vl_types.all;
entity keyMatrix_test is
end keyMatrix_test;
