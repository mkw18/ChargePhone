library verilog;
use verilog.vl_types.all;
entity mechine_test is
end mechine_test;
