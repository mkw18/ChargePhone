library verilog;
use verilog.vl_types.all;
entity setNum_vlg_vec_tst is
end setNum_vlg_vec_tst;
