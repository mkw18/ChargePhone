library verilog;
use verilog.vl_types.all;
entity scan_vlg_vec_tst is
end scan_vlg_vec_tst;
